`timescale 1ns/1ps

module CRC_tb;

/////////////////////////////////////////////////////////
///////////////////// Parameters ////////////////////////
/////////////////////////////////////////////////////////

parameter period = 100;
parameter DWIDTH = 8;
parameter DDEPTH = 10;

/////////////////////////////////////////////////////////
///////////////////// Declaratios ///////////////////////
/////////////////////////////////////////////////////////

reg     data_tb;
reg     active_tb;
reg     clk_tb;
reg     rst_tb;
wire    crc_tb;
wire    valid_tb;

/////////////////////////////////////////////////////////
//////////////////////// Vars ///////////////////////////
/////////////////////////////////////////////////////////

integer i=0;
reg     [DWIDTH-1:0] gener_out;

/////////////////////////////////////////////////////////
///////////////////// memories //////////////////////////
/////////////////////////////////////////////////////////

reg     [DWIDTH-1:0]     mem     [DDEPTH-1:0];
reg     [DWIDTH-1:0]     rus     [DDEPTH-1 :0];

/////////////////////////////////////////////////////////
///////////////////// Instantiation /////////////////////
/////////////////////////////////////////////////////////

CRC DUT(data_tb, active_tb, clk_tb, rst_tb, crc_tb, valid_tb);

/////////////////////////////////////////////////////////
///////////////////// Clock generation //////////////////
/////////////////////////////////////////////////////////

always #(0.5 * period) clk_tb = ~clk_tb;

/////////////////////////////////////////////////////////
///////////////////// Initial Block /////////////////////
/////////////////////////////////////////////////////////

initial begin
    //System functions.
    $dumpfile("LFSR_DUMP.vcd") ;       
    $dumpvars; 

    //Read files.
    $readmemh("DATA_h.txt",mem);
    $readmemh("Expec_Out_h.txt",rus);
    
    //initialization.
    init;

    for(i=0; i<10; i=i+1)
    begin
        do_oper(mem[i]);    //do the operation for each byte in mem.
        check(i);           //Check the output.
    end

    #(20 * period)
    $stop;
end

/////////////////////////////////////////////////////////
///////////////////// Tasks /////////////////////////////
/////////////////////////////////////////////////////////

/////////////// Signals Initialization //////////////////
task init;
begin
    clk_tb = 'b0;
    rst_tb = 'b0;
    active_tb = 'b0;
end
endtask

//////////////////////// Reset /////////////////////////
task reset;
begin
    rst_tb = 'b1;
    #period;
    rst_tb = 'b0;
end
endtask

////////////////// Do LFSR Operation ////////////////////
task do_oper;
input [DWIDTH-1:0] byte;
integer x;
begin
    reset;
    active_tb = 'b1;

    for(x=0; x<DWIDTH; x=x+1)
    begin
        data_tb = byte[x];
        #period;
    end
    get_out;
end
endtask

////////////// Store the output of the CRC //////////////
task get_out;
integer j;
begin
    active_tb = 'b0;
    @(posedge valid_tb)
    for(j=0; j<DWIDTH; j=j+1)
    begin
        #period gener_out[j] = crc_tb;
    end    
end
endtask 

////////////////// Check Out Response  //////////////////
task check;
input integer z;
begin
    if(gener_out == rus[z])
        $display("test number %0d is passed",i);
    else
        $display("test number %0d is failed",i);
end
endtask


endmodule